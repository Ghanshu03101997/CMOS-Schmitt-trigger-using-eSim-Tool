* C:\Users\lenovo\eSim-Workspace\Schmitt_Trigger\Schmitt_Trigger.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 09-Mar-22 9:19:44 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M3  Net-_M3-Pad1_ in Net-_M3-Pad3_ Net-_M3-Pad1_ eSim_MOS_P		
M4  Net-_M3-Pad3_ in out Net-_M3-Pad3_ eSim_MOS_P		
M1  out in Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
M2  Net-_M1-Pad3_ in Net-_M2-Pad3_ Net-_M2-Pad3_ eSim_MOS_N		
M6  Net-_M6-Pad1_ out Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
M5  Net-_M3-Pad3_ out GND Net-_M3-Pad3_ eSim_MOS_P		
v2  Net-_M3-Pad1_ GND 1.8		
v3  Net-_M6-Pad1_ Net-_M2-Pad3_ 1.8		
U2  out plot_v1		
U1  in plot_v1		
v1  in GND 1.8		

.end
